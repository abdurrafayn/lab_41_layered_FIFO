always_ff @( edge clk ) begin : slowclock
    
end